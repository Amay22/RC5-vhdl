LIBRARY	IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;


PACKAGE rc5_pkg IS
TYPE ROM1 IS ARRAY(0 TO 25) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
END rc5_pkg;
